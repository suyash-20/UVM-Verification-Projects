package seq_package;


import uvm_pkg::*;

`include "uvm_macros.svh"

	`include "trans_xtn.sv"
	`include "seq_agent_config.sv"

	`include "seq_env_config.sv"


	`include "driver_callback.sv"  //CALLBACK LOGIC
	`include "custom_callback.sv"  //CALLBACK LOGIC

	`include "seq_driver.sv"
	`include "seq_monitor.sv"
	`include "seq_sequencer.sv"
	`include "seq_agent.sv"
	`include "seq_agt_top.sv"
	`include "seq_sequence.sv"


	`include "virtual_sequencer.sv"
	`include "virtual_sequence.sv"
	`include "seq_scoreboard.sv"

	
	`include "seq_tb.sv"
	`include "seq_test.sv"

endpackage

